module _32bit_mux_2x1 (R, S, I0, I1);
input S;
input [31:0] I0, I1;
output [31:0] R;

mux_2x1  mux0(R[0], S, I0[0], I1[0]),
			mux1(R[1], S, I0[1], I1[1]),
			mux2(R[2], S, I0[2], I1[2]),
			mux3(R[3], S, I0[3], I1[3]),
			mux4(R[4], S, I0[4], I1[4]),
			mux5(R[5], S, I0[5], I1[5]),
			mux6(R[6], S, I0[6], I1[6]),
			mux7(R[7], S, I0[7], I1[7]),
			mux8(R[8], S, I0[8], I1[8]),
			mux9(R[9], S, I0[9], I1[9]),
			mux10(R[10], S, I0[10], I1[10]),
			mux11(R[11], S, I0[11], I1[11]),
			mux12(R[12], S, I0[12], I1[12]),
			mux13(R[13], S, I0[13], I1[13]),
			mux14(R[14], S, I0[14], I1[14]),
			mux15(R[15], S, I0[15], I1[15]),
			mux16(R[16], S, I0[16], I1[16]),
			mux17(R[17], S, I0[17], I1[17]),
			mux18(R[18], S, I0[18], I1[18]),
			mux19(R[19], S, I0[19], I1[19]),
			mux20(R[20], S, I0[20], I1[20]),
			mux21(R[21], S, I0[21], I1[21]),
			mux22(R[22], S, I0[22], I1[22]),
			mux23(R[23], S, I0[23], I1[23]),
			mux24(R[24], S, I0[24], I1[24]),
			mux25(R[25], S, I0[25], I1[25]),
			mux26(R[26], S, I0[26], I1[26]),
			mux27(R[27], S, I0[27], I1[27]),
			mux28(R[28], S, I0[28], I1[28]),
			mux29(R[29], S, I0[29], I1[29]),
			mux30(R[30], S, I0[30], I1[30]),
			mux31(R[31], S, I0[31], I1[31]);

endmodule
