module sign_extend(R, I);
input [5:0] I;
output [31:0] R;

mux_2x1 mux31(R[31], I[5], 1'b0, 1'b1),
		  mux30(R[30], I[5], 1'b0, 1'b1),
		  mux29(R[29], I[5], 1'b0, 1'b1),
		  mux28(R[28], I[5], 1'b0, 1'b1),
	 	  mux27(R[27], I[5], 1'b0, 1'b1),
		  mux26(R[26], I[5], 1'b0, 1'b1),
		  mux25(R[25], I[5], 1'b0, 1'b1),
		  mux24(R[24], I[5], 1'b0, 1'b1),
		  mux23(R[23], I[5], 1'b0, 1'b1),
		  mux22(R[22], I[5], 1'b0, 1'b1),
		  mux21(R[21], I[5], 1'b0, 1'b1),
		  mux20(R[20], I[5], 1'b0, 1'b1),
		  mux19(R[19], I[5], 1'b0, 1'b1),
		  mux18(R[18], I[5], 1'b0, 1'b1),
		  mux17(R[17], I[5], 1'b0, 1'b1),
		  mux16(R[16], I[5], 1'b0, 1'b1),
		  mux15(R[15], I[5], 1'b0, 1'b1),
		  mux14(R[14], I[5], 1'b0, 1'b1),
		  mux13(R[13], I[5], 1'b0, 1'b1),
		  mux12(R[12], I[5], 1'b0, 1'b1),
		  mux11(R[11], I[5], 1'b0, 1'b1),
		  mux10(R[10], I[5], 1'b0, 1'b1),
		  mux9(R[9], I[5], 1'b0, 1'b1),
		  mux8(R[8], I[5], 1'b0, 1'b1),
		  mux7(R[7], I[5], 1'b0, 1'b1),
		  mux6(R[6], I[5], 1'b0, 1'b1);
		  
or or5(R[5], I[5], 1'b0),
	or4(R[4], I[4], 1'b0),
	or3(R[3], I[3], 1'b0),
	or2(R[2], I[2], 1'b0),
	or1(R[1], I[1], 1'b0),
	or0(R[0], I[0], 1'b0);

endmodule
