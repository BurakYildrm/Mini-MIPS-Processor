module _32bit_mux_8x1 (R, S2, S1, S0, I0, I1, I2, I3, I4, I5, I6, I7);
input S2, S1, S0;
input [31:0] I0, I1, I2, I3, I4, I5, I6, I7;
output [31:0] R;

mux_8x1  mux0(R[0], S2, S1, S0, I0[0], I1[0], I2[0], I3[0], I4[0], I5[0], I6[0], I7[0]),
         mux1(R[1], S2, S1, S0, I0[1], I1[1], I2[1], I3[1], I4[1], I5[1], I6[1], I7[1]),
         mux2(R[2], S2, S1, S0, I0[2], I1[2], I2[2], I3[2], I4[2], I5[2], I6[2], I7[2]),
         mux3(R[3], S2, S1, S0, I0[3], I1[3], I2[3], I3[3], I4[3], I5[3], I6[3], I7[3]),
         mux4(R[4], S2, S1, S0, I0[4], I1[4], I2[4], I3[4], I4[4], I5[4], I6[4], I7[4]),
         mux5(R[5], S2, S1, S0, I0[5], I1[5], I2[5], I3[5], I4[5], I5[5], I6[5], I7[5]),
         mux6(R[6], S2, S1, S0, I0[6], I1[6], I2[6], I3[6], I4[6], I5[6], I6[6], I7[6]),
         mux7(R[7], S2, S1, S0, I0[7], I1[7], I2[7], I3[7], I4[7], I5[7], I6[7], I7[7]),
         mux8(R[8], S2, S1, S0, I0[8], I1[8], I2[8], I3[8], I4[8], I5[8], I6[8], I7[8]),
         mux9(R[9], S2, S1, S0, I0[9], I1[9], I2[9], I3[9], I4[9], I5[9], I6[9], I7[9]),
         mux10(R[10], S2, S1, S0, I0[10], I1[10], I2[10], I3[10], I4[10], I5[10], I6[10], I7[10]),
         mux11(R[11], S2, S1, S0, I0[11], I1[11], I2[11], I3[11], I4[11], I5[11], I6[11], I7[11]),
         mux12(R[12], S2, S1, S0, I0[12], I1[12], I2[12], I3[12], I4[12], I5[12], I6[12], I7[12]),
         mux13(R[13], S2, S1, S0, I0[13], I1[13], I2[13], I3[13], I4[13], I5[13], I6[13], I7[13]),
         mux14(R[14], S2, S1, S0, I0[14], I1[14], I2[14], I3[14], I4[14], I5[14], I6[14], I7[14]),
         mux15(R[15], S2, S1, S0, I0[15], I1[15], I2[15], I3[15], I4[15], I5[15], I6[15], I7[15]),
         mux16(R[16], S2, S1, S0, I0[16], I1[16], I2[16], I3[16], I4[16], I5[16], I6[16], I7[16]),
         mux17(R[17], S2, S1, S0, I0[17], I1[17], I2[17], I3[17], I4[17], I5[17], I6[17], I7[17]),
         mux18(R[18], S2, S1, S0, I0[18], I1[18], I2[18], I3[18], I4[18], I5[18], I6[18], I7[18]),
         mux19(R[19], S2, S1, S0, I0[19], I1[19], I2[19], I3[19], I4[19], I5[19], I6[19], I7[19]),
         mux20(R[20], S2, S1, S0, I0[20], I1[20], I2[20], I3[20], I4[20], I5[20], I6[20], I7[20]),
         mux21(R[21], S2, S1, S0, I0[21], I1[21], I2[21], I3[21], I4[21], I5[21], I6[21], I7[21]),
         mux22(R[22], S2, S1, S0, I0[22], I1[22], I2[22], I3[22], I4[22], I5[22], I6[22], I7[22]),
         mux23(R[23], S2, S1, S0, I0[23], I1[23], I2[23], I3[23], I4[23], I5[23], I6[23], I7[23]),
         mux24(R[24], S2, S1, S0, I0[24], I1[24], I2[24], I3[24], I4[24], I5[24], I6[24], I7[24]),
         mux25(R[25], S2, S1, S0, I0[25], I1[25], I2[25], I3[25], I4[25], I5[25], I6[25], I7[25]),
         mux26(R[26], S2, S1, S0, I0[26], I1[26], I2[26], I3[26], I4[26], I5[26], I6[26], I7[26]),
         mux27(R[27], S2, S1, S0, I0[27], I1[27], I2[27], I3[27], I4[27], I5[27], I6[27], I7[27]),
         mux28(R[28], S2, S1, S0, I0[28], I1[28], I2[28], I3[28], I4[28], I5[28], I6[28], I7[28]),
         mux29(R[29], S2, S1, S0, I0[29], I1[29], I2[29], I3[29], I4[29], I5[29], I6[29], I7[29]),
         mux30(R[30], S2, S1, S0, I0[30], I1[30], I2[30], I3[30], I4[30], I5[30], I6[30], I7[30]),
         mux31(R[31], S2, S1, S0, I0[31], I1[31], I2[31], I3[31], I4[31], I5[31], I6[31], I7[31]);

endmodule
